module rom #(
    parameter   ADD_WIDTH = 8,
                DATA_WIDTH = 8
)(
    input logic clk,
    input logic [ADD_WIDTH-1:0] addr,
    input logic [ADD_WIDTH-1:0] addr2,
    output logic [DATA_WIDTH-1:0] dout,
    output logic [DATA_WIDTH-1:0] dout2

);

logic [DATA_WIDTH-1:0] rom_array [2**ADD_WIDTH-1:0];

initial begin
    $display("Loading rom.");
    $readmemh("sinerom.mem",rom_array);

end;

always_ff @ (posedge clk) 
begin
    dout <= rom_array [addr];
    dout2 <= rom_array [addr2];
end
endmodule
